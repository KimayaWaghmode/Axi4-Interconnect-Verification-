These are the verification files for AXI4 Interconnect Verification
