Adding the design files for AXI4 Interconnect Verification
