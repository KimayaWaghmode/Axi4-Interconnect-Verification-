Design files for AXI4 Interconnect Verification
